`timescale 1ns/1ps

module tb_hpu_cmp_node ();


endmodule