module gcu_top (


    input logic clk,
    input logic rstn
);
    
endmodule