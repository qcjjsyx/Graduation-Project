`timescale 1ns/1ps

module tb_hpu_core_tree ();


endmodule